module hvif
